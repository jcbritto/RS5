/*!\file testbench.sv
 * RS5 VERSION - 1.1.0 - Pipeline Simplified and Core Renamed
 *
 * Distribution:  October 2023
 *
 * Willian Nunes    <willian.nunes@edu.pucrs.br>
 * Angelo Dal Zotto <angelo.dalzotto@edu.pucrs.br>
 * Marcos Sartori   <marcos.sartori@acad.pucrs.br>
 * Ney Calazans     <ney.calazans@ufsc.br>
 * Fernando Moraes  <fernando.moraes@pucrs.br>
 * GAPH - Hardware Design Support Group
 * PUCRS - Pontifical Catholic University of Rio Grande do Sul <https://pucrs.br/>
 *
 * \brief
 * Testbench for RS5 simulation.
 *
 * \detailed
 * Testbench for RS5 simulation.de
 */

`include "../rtl/RS5_pkg.sv"

//////////////////////////////////////////////////////////////////////////////
// CPU TESTBENCH
//////////////////////////////////////////////////////////////////////////////

module testbench
    import RS5_pkg::*;
(
);
    timeunit 1ns; timeprecision 1ns;

//////////////////////////////////////////////////////////////////////////////
// PARAMETERS FOR CORE INSTANTIATION
//////////////////////////////////////////////////////////////////////////////

    localparam mul_e         MULEXT          = MUL_M;
    localparam atomic_e      AMOEXT          = AMO_A;
    localparam bit           COMPRESSED      = 1'b1;
    localparam bit           USE_XOSVM       = 1'b0;
    localparam bit           USE_ZKNE        = 1'b1;
    localparam bit           USE_ZICOND      = 1'b1;
    localparam bit           USE_ZCB         = 1'b1;
    localparam bit           VEnable         = 1'b0;
    localparam int           VLEN            = 256;
    localparam int           LLEN            = 32;
    localparam bit           USE_HPMCOUNTER  = 1'b1;
    localparam bit           BRANCHPRED      = 1'b1;
    localparam bit           FORWARDING      = 1'b1;

`ifndef SYNTH
    localparam bit           PROFILING       = 1'b1;
    localparam bit           DEBUG           = 1'b0;
`endif
    localparam string        PROFILING_FILE  = "./results/Report.txt";
    localparam string        OUTPUT_FILE     = "./results/Output.txt";

    localparam int           MEM_WIDTH       = 65_536;
    localparam string        BIN_FILE        = "./test_debug_c.bin";

    localparam int           i_cnt = 1;

///////////////////////////////////////// Clock generator //////////////////////////////

    logic        clk=1;

    always begin
        #5.0 clk <= 0;
        #5.0 clk <= 1;
    end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// RESET CPU ////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

    logic reset_n;

    // Basic debug - count any memory write operation
    integer write_count = 0;
    always_ff @(posedge clk) begin
        if (mem_write_enable != '0) begin
            write_count <= write_count + 1;
            $display("# %0t Memory Write %0d: addr=0x%08X, data=0x%08X, enable=0x%X", 
                     $time, write_count, mem_address, mem_data_write, mem_write_enable);
        end
        
        // Debug ADD_PLUGIN instruction detection
        if (dut.decoder1.instruction_i[6:0] == 7'b0001011) begin
            $display("# %0t CUSTOM-0 Instruction: 0x%08X", $time, dut.decoder1.instruction_i);
        end
        if (dut.execute1.instruction_operation_i == ADD_PLUGIN) begin
            $display("# %d ADD_PLUGIN Operation Detected!", $time);
            $display("# %d   Instruction: 0x%08x", $time, dut.execute1.instruction_i);
            $display("# %d   rs1=x%0d, rs2=x%0d, rd=x%0d", $time, 
                     dut.execute1.instruction_i[19:15],
                     dut.execute1.instruction_i[24:20], 
                     dut.execute1.instruction_i[11:7]);
            $display("# %d   op_a_value=0x%08x, op_b_value=0x%08x", $time,
                     dut.execute1.rs1_data_i,
                     dut.execute1.rs2_data_i);
        end
        
        // Debug plugin execution in execute stage
        if (dut.execute1.plugin_enable) begin
            $display("# %0t Plugin Enable: start=%b, busy=%b, done=%b, op_a=0x%08X, op_b=0x%08X, result=0x%08X", 
                     $time, dut.execute1.plugin_start, dut.execute1.plugin_busy, dut.execute1.plugin_done,
                     dut.execute1.rs1_data_i, dut.execute1.rs2_data_i, dut.execute1.plugin_result);
        end
    end

    initial begin
        reset_n = 0;                                          // RESET for CPU initialization

        #100 reset_n = 1;                                     // Hold state for 100 ns
        
        // Timeout para evitar simulação infinita
        #500000 begin
            $display("\n# %0t TIMEOUT - ENDING SIMULATION", $time);
            $finish;
        end
    end

//////////////////////////////////////////////////////////////////////////////
// TB SIGNALS
//////////////////////////////////////////////////////////////////////////////

    /* Number of used bits is defined by the memory size */
    /* verilator lint_off UNUSEDSIGNAL */
    logic [31:0]            instruction_address;
    /* verilator lint_on UNUSEDSIGNAL */

    /* RTC is 64 bits but the bus is 32 bits */
    /* verilator lint_off UNUSEDSIGNAL */
    logic [63:0]            data_rtc;
    /* verilator lint_on UNUSEDSIGNAL */

    logic                   interrupt_ack;
    logic [63:0]            mtime;
    logic [31:0]            instruction;
    logic                   enable_ram, enable_rtc, enable_plic, enable_tb, enable_plugin;
    logic                   mem_operation_enable;
    logic [31:0]            mem_address, mem_data_read, mem_data_write;
    logic [3:0]             mem_write_enable;
    byte                    char;
    logic [31:0]            data_ram, data_plic, data_tb, data_plugin;
    logic                   enable_tb_r, enable_rtc_r, enable_plic_r, enable_plugin_r;
    logic                   mti, mei;

//////////////////////////////////////////////////////////////////////////////
// Control
//////////////////////////////////////////////////////////////////////////////

    always_comb begin
        if (mem_operation_enable) begin
            if (mem_address[31:28] < 4'h1) begin
                enable_ram    = 1'b1;
                enable_plugin = 1'b0;
                enable_rtc    = 1'b0;
                enable_plic   = 1'b0;
                enable_tb     = 1'b0;
            end
            else if (mem_address[31:28] < 4'h2) begin
                enable_ram    = 1'b0;
                enable_plugin = 1'b1;
                enable_rtc    = 1'b0;
                enable_plic   = 1'b0;
                enable_tb     = 1'b0;
            end
            else if (mem_address[31:28] < 4'h3) begin
                enable_ram    = 1'b0;
                enable_plugin = 1'b0;
                enable_rtc    = 1'b1;
                enable_plic   = 1'b0;
                enable_tb     = 1'b0;
            end
            else if (mem_address[31:28] < 4'h8) begin
                enable_ram    = 1'b0;
                enable_plugin = 1'b0;
                enable_rtc    = 1'b0;
                enable_plic   = 1'b1;
                enable_tb     = 1'b0;
            end
            else begin
                enable_ram    = 1'b0;
                enable_plugin = 1'b0;
                enable_rtc    = 1'b0;
                enable_plic   = 1'b0;
                enable_tb     = 1'b1;
            end
        end
        else begin
            enable_ram    = 1'b0;
            enable_plugin = 1'b0;
            enable_rtc    = 1'b0;
            enable_plic   = 1'b0;
            enable_tb     = 1'b0;
        end
    end

    always_ff @(posedge clk) begin
        enable_tb_r     <= enable_tb;
        enable_rtc_r    <= enable_rtc;
        enable_plic_r   <= enable_plic;
        enable_plugin_r <= enable_plugin;
    end

    always_comb begin
        if (enable_tb_r) begin
            mem_data_read = data_tb;
        end
        else if (enable_rtc_r) begin
            mem_data_read = data_rtc[31:0];
        end
        else if (enable_plic_r) begin
            mem_data_read = data_plic;
        end
        else if (enable_plugin_r) begin
            mem_data_read = data_plugin;
        end
        else begin
            mem_data_read = data_ram;
        end
    end

//////////////////////////////////////////////////////////////////////////////
// CPU
//////////////////////////////////////////////////////////////////////////////

    RS5 #(
    `ifndef SYNTH
	    .DEBUG          (DEBUG          ),
	    .PROFILING      (PROFILING      ),
        .PROFILING_FILE (PROFILING_FILE ),
    `endif
        .Environment     (ASIC          ),
        .MULEXT          (MULEXT        ),
        .AMOEXT          (AMOEXT        ),
        .COMPRESSED      (COMPRESSED    ),
        .VEnable         (VEnable       ),
        .VLEN            (VLEN          ),
        .LLEN            (LLEN          ),
        .XOSVMEnable     (USE_XOSVM     ),
        .ZKNEEnable      (USE_ZKNE      ),
        .ZICONDEnable    (USE_ZICOND    ),
        .ZCBEnable       (USE_ZCB       ),
        .HPMCOUNTEREnable(USE_HPMCOUNTER),
        .BRANCHPRED      (BRANCHPRED    ),
        .FORWARDING      (FORWARDING    )
    ) dut (
        .clk                    (clk),
        .reset_n                (reset_n),
        .sys_reset_i            (1'b0),
        .stall                  (1'b0),
        .instruction_i          (instruction),
        .mem_data_i             (mem_data_read),
        .mtime_i                (mtime),
        .tip_i                  (mti),
        .eip_i                  (mei),
        .instruction_address_o  (instruction_address),
        .mem_operation_enable_o (mem_operation_enable),
        .mem_write_enable_o     (mem_write_enable),
        .mem_address_o          (mem_address),
        .mem_data_o             (mem_data_write),
        .interrupt_ack_o        (interrupt_ack)
    );

//////////////////////////////////////////////////////////////////////////////
// RAM
//////////////////////////////////////////////////////////////////////////////

    RAM_mem #(
    `ifndef SYNTH
        .DEBUG     (DEBUG     ),
        .DEBUG_PATH("./debug/"),
    `endif
        .MEM_WIDTH(MEM_WIDTH  ),
        .BIN_FILE (BIN_FILE   )
    ) RAM_MEM (
        .clk        (clk),

        .enA_i      (1'b1),
        .weA_i      (4'h0),
        .addrA_i    (instruction_address[($clog2(MEM_WIDTH) - 1):0]),
        .dataA_i    (32'h00000000),
        .dataA_o    (instruction),

        .enB_i      (enable_ram),
        .weB_i      (mem_write_enable),
        .addrB_i    (mem_address[($clog2(MEM_WIDTH) - 1):0]),
        .dataB_i    (mem_data_write),
        .dataB_o    (data_ram)
    );

//////////////////////////////////////////////////////////////////////////////
// PLIC
//////////////////////////////////////////////////////////////////////////////

    /* Bits depending on connected peripherals */
    /* verilator lint_off UNUSED */
    logic [i_cnt:1] iack_periph;
    /* verilator lint_on UNUSED */

    plic #(
        .i_cnt(i_cnt)
    ) plic1 (
        .clk     (clk),
        .reset_n (reset_n),
        .en_i    (enable_plic),
        .we_i    (mem_write_enable),
        .addr_i  (mem_address[23:0]),
        .data_i  (mem_data_write),
        .data_o  (data_plic),
        .irq_i   ('0),
        .iack_i  (interrupt_ack),
        .iack_o  (iack_periph),
        .irq_o   (mei)
    );

//////////////////////////////////////////////////////////////////////////////
// RTC
//////////////////////////////////////////////////////////////////////////////

    rtc rtc(
        .clk        (clk),
        .reset_n    (reset_n),
        .en_i       (enable_rtc),
        .addr_i     (mem_address[3:0]),
        .we_i       ({4'h0, mem_write_enable}),
        .data_i     ({32'h0, mem_data_write}),
        .data_o     (data_rtc),
        .mti_o      (mti),
        .mtime_o    (mtime)
    );

//////////////////////////////////////////////////////////////////////////////
// PLUGIN
//////////////////////////////////////////////////////////////////////////////

    plugin_memory_interface plugin_mem_if(
        .clk      (clk),
        .reset_n  (reset_n),
        .enable_i (enable_plugin),
        .we_i     (mem_write_enable),
        .addr_i   (mem_address),
        .data_i   (mem_data_write),
        .data_o   (data_plugin)
    );

//////////////////////////////////////////////////////////////////////////////
// Memory Mapped regs
//////////////////////////////////////////////////////////////////////////////
    int fd;
    initial begin
        fd = $fopen(OUTPUT_FILE,"w");
    end

    always_ff @(posedge clk) begin
        if (enable_tb) begin
            // OUTPUT REG
            if ((mem_address == 32'h80004000 || mem_address == 32'h80001000) && mem_write_enable != '0) begin
                char <= mem_data_write[7:0];
                $write("%c",char);
                if (char != 8'h00)
                    $fwrite(fd,"%c",char);
                $fflush();
            end
            else if (mem_address == 32'h80002000 && mem_write_enable != '0) begin
                $write(    "%0d\n",mem_data_write);
                $fwrite(fd,"%0d\n",mem_data_write);
                $fflush();
            end
            // ADD_PLUGIN TEST DEBUG
            else if ((mem_address >= 32'h00001000 && mem_address < 32'h00001010) && mem_write_enable != '0) begin
                $display("# %0t ADD_PLUGIN Test: Writing 0x%08X to address 0x%08X", $time, mem_data_write, mem_address);
            end
            // END REG
            if (mem_address == 32'h80000000 && mem_write_enable != '0) begin
                $display(    "\n# %0t END OF SIMULATION",$time);
                $fdisplay(fd,"\n# %0t END OF SIMULATION",$time);
                $finish;
            end
        end
        else begin
            data_tb <= '0;
        end
    end

endmodule
